module TS_STATE_MACHINE(
	
	input SYS_CLOCK			,
	input SYS_RESET			,

	input TS_CLOCK_IN			,
	input TS_RESET				,
	
	input PASS					,
	input PLAY					,
	input REC					,
	
	input			TS_VALID_IN	,
	input			TS_SYNC_IN	,
	input	 [7:0]TS_DATA_IN	,
	
	output		TS_VALID_OUT,
	output		TS_SYNC_OUT	,
	output [7:0]TS_DATA_OUT	,
	
	output 		TS_CLOCK_OUT,
	
	output reg [1:0] STATE
);

wire			B_VALID	;
wire			B_SYNC	;
wire	[7:0]	B_DATA	;

BUFFER_IP #(
	.WIDTH		(10)
	)
	TS_BUFFER_IP(
	.CLOCK		(TS_CLOCK_IN										),
	.RESET		(TS_RESET											),
	.DATA_IN		({TS_VALID_IN, TS_SYNC_IN, TS_DATA_IN}		),
	.DATA_OUT	({B_VALID, B_SYNC, B_DATA}						)
);

reg			TEMP_VALID	;
reg			TEMP_SYNC	;
reg	[7:0]	TEMP_DATA	;

localparam PASSTHROUGH	= 2'b00;
localparam RECORD			= 2'b01;
localparam REPLAY			= 2'b10;

always @(posedge SYS_CLOCK or posedge SYS_RESET)	begin

	if(SYS_RESET)	begin
	
		STATE <= PASSTHROUGH;
	end
	else	begin
	
		case(STATE)
		
			PASSTHROUGH:	begin
				
				if(PLAY || REC)	begin
				
					if(PLAY	)	STATE <= REPLAY;
					if(REC	)	STATE <= RECORD;
				end
				else	begin
				
					STATE <= PASSTHROUGH;
				end
				
				TEMP_VALID	= B_VALID	;
				TEMP_SYNC	= B_SYNC		;
				TEMP_DATA	= B_DATA		;
			end
			
			RECORD:	begin
			
				STATE <= (PASS	)? PASSTHROUGH : RECORD;
				
				TEMP_VALID	= B_VALID	;
				TEMP_SYNC	= B_SYNC		;
				TEMP_DATA	= B_DATA		;
			end
			
			REPLAY:	begin
			
				STATE <= (PASS	)? PASSTHROUGH : REPLAY;
			end
		endcase
	end
end

BUFFER_COMB #(
	.WIDTH		(10)
	)
	TS_BUFFER_OP(
	.CLOCK		(TS_CLOCK_IN										),
	.RESET		(TS_RESET											),
	.DATA_IN		({TEMP_VALID, TEMP_SYNC, TEMP_DATA}			),
	.DATA_OUT	({TS_VALID_OUT, TS_SYNC_OUT, TS_DATA_OUT}	)
);

assign	TS_CLOCK_OUT	= TS_CLOCK_IN	;



//BUFFER_COMB #(
//	.WIDTH		(10)
//	)
//	TS_BUFFER(
//	.CLOCK		(TS_CLOCK_IN										),
//	.RESET		(TS_RESET											),
//	.DATA_IN		({TS_VALID_IN, TS_SYNC_IN, TS_DATA_IN}		),
//	.DATA_OUT	({TS_VALID_OUT, TS_SYNC_OUT, TS_DATA_OUT}	)
//);

//assign TS_VALID_OUT	= TEMP_VALID;
//assign TS_SYNC_OUT	= TEMP_SYNC	;
//assign TS_DATA_OUT	= TEMP_DATA	;


//
//assign	TS_VALID_OUT	= TS_VALID_IN	;
//assign	TS_SYNC_OUT		= TS_SYNC_IN	;
//
//assign	TS_DATA_OUT		= TS_DATA_IN	;

endmodule
