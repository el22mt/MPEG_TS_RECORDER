module TS_BUFFER #(
	parameter WIDTH = 10
	)(
	input							CLOCK		,
	input							RESET		,
	input		  [WIDTH-1 : 0]DATA_IN	,
	
	output reg [WIDTH-1 : 0]DATA_OUT
);

always @(posedge CLOCK or posedge RESET)	begin

	if(RESET)	begin
	
		DATA_OUT <= {WIDTH{1'b0}}	;
	end
	else	begin
	
		DATA_OUT <= DATA_IN			;
	end
end
endmodule
